#single upper case letter are usually initials
A
B
C
D
E
F
G
H
I
J
K
L
M
N
O
P
Q
R
S
T
U
V
W
X
Y
Z
#misc abbreviations
AB
G
VG
dvs
etc
from
iaf
jfr
kl
kr
mao
mfl
mm
osv
pga
tex
tom
vs
